// You need to generate this component correctly

module dmem(addr,clk,data,wren,q);

input clk,wren;
input [11:0] addr;
input [31:0] data;
output [31:0] q;

endmodule
