// You need to generate this component correctly
module imem(addr,clk,q);

input clk;
input [11:0] addr;
output reg[31:0] q;

always @(posedge clk) begin
	
end

endmodule
